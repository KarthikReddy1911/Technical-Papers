module full_adder(input a,b,c,output sum,cout);
 logic a,b,c;
 logic sum,cout;
 assign {cout,sum}=a+b+c;
endmodule
//thank you
//jaswanth 
